CIRCUIT example
*
* IC Technology: CMOS 0.12�m - 6 Metal
*
VDD 1 0 DC 1.20
*
* List of nodes
*
* MOS devices
*
*
*
* Transient analysis
*
.TEMP 27.0
.TRAN 0.1N 5.00N
* (Pspice)
.PROBE
.END
